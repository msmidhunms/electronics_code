library IEEE;
use IEEE.std_logic.all;
