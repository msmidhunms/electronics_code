library IEEE;
use IEEE.std_logic.all;
entity simple is
      port(a,b : in std_logic; c: out std_logic);
end entity simple

architecture behaviour of simple is
begin

end behaviour
